module my_and(input in_a,
              input in_b,
              output out);
    
    assign out = in_a & in_b;
    // and and_1(out, in_a, in_b);  
  
endmodule 
